library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity comb_logic is
	port(	i_a
		i_b
		O-c 
