library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity reg is
   port (clk : in std_logic := '0';
         reset : in std_logic := '0';
         
         i_d : in std_logic := '0';
         
         o_q : out std_logic := '0');
end reg;



architecture rtl of reg is
  
--signal declaration
  
  
begin

--synchronous process
   process (clk) is
   begin
      if rising_edge(clk) then  
        if (reset='1') then   
            o_q <= '0';
         else
            o_q <= i_d; 
      	end if;
      end if;
   end process;



end rtl;
